// Instanciamos en el core y conectamos los registros de segmentación. Podrán ser descritos directamente en el módulo top mediante bloques procedimentales always.


